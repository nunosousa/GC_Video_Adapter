-- file: gc_dv_top_level.vhd

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity gc_dv_top_level is
	port(

	);
	
end entity;

architecture behav of gc_dv_top_level is
	
begin

end behav;

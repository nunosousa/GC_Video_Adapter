-- file: gc_dv_decode_tb.vhd
